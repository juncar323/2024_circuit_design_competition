`timescale 1ns / 1ps

module layer_3 #(
DATA_WIDTH = 32
)(
    input logic [DATA_WIDTH-1:0] data0,   // 채널 0의 입력 데이터
    input logic [DATA_WIDTH-1:0] data1,   // 채널 1의 입력 데이터
    input logic [DATA_WIDTH-1:0] data2,   // 채널 2의 입력 데이터
    input logic [DATA_WIDTH-1:0] data3,   // 채널 3의 입력 데이터
    input logic [DATA_WIDTH-1:0] data4,   // 채널 4의 입력 데이터
    input logic [DATA_WIDTH-1:0] data5,   // 채널 5의 입력 데이터
    input logic [DATA_WIDTH-1:0] data6,   // 채널 6의 입력 데이터
    input logic [DATA_WIDTH-1:0] data7,   // 채널 7의 입력 데이터
    input logic [DATA_WIDTH-1:0] data8,   // 채널 8의 입력 데이터
    input logic [DATA_WIDTH-1:0] data9,   // 채널 9의 입력 데이터
    input logic [DATA_WIDTH-1:0] data10,  // 채널 10의 입력 데이터
    input logic [DATA_WIDTH-1:0] data11,  // 채널 11의 입력 데이터
    input logic [DATA_WIDTH-1:0] data12,  // 채널 12의 입력 데이터
    input logic [DATA_WIDTH-1:0] data13,  // 채널 13의 입력 데이터
    input logic [DATA_WIDTH-1:0] data14,  // 채널 14의 입력 데이터
    input logic [DATA_WIDTH-1:0] data15,  // 채널 15의 입력 데이터
    input logic [DATA_WIDTH-1:0] data16,  // 채널 16의 입력 데이터
    input logic [DATA_WIDTH-1:0] data17,  // 채널 17의 입력 데이터
    input logic [DATA_WIDTH-1:0] data18,  // 채널 18의 입력 데이터
    input logic [DATA_WIDTH-1:0] data19,  // 채널 19의 입력 데이터
    input logic [DATA_WIDTH-1:0] data20,  // 채널 20의 입력 데이터
    input logic [DATA_WIDTH-1:0] data21,  // 채널 21의 입력 데이터
    input logic [DATA_WIDTH-1:0] data22,  // 채널 22의 입력 데이터
    input logic [DATA_WIDTH-1:0] data23,  // 채널 23의 입력 데이터
    input logic [DATA_WIDTH-1:0] data24,  // 채널 24의 입력 데이터
    input logic [DATA_WIDTH-1:0] data25,  // 채널 25의 입력 데이터
    input logic [DATA_WIDTH-1:0] data26,  // 채널 26의 입력 데이터
    input logic [DATA_WIDTH-1:0] data27,  // 채널 27의 입력 데이터
    input logic [DATA_WIDTH-1:0] data28,  // 채널 28의 입력 데이터
    input logic [DATA_WIDTH-1:0] data29,  // 채널 29의 입력 데이터
    input logic [DATA_WIDTH-1:0] data30,  // 채널 30의 입력 데이터
    input logic [DATA_WIDTH-1:0] data31,
    input logic [DATA_WIDTH-1:0] data32,
    input logic [DATA_WIDTH-1:0] data33,
    input logic [DATA_WIDTH-1:0] data34,
    input logic [DATA_WIDTH-1:0] data35,
    input logic [DATA_WIDTH-1:0] data36,
    input logic [DATA_WIDTH-1:0] data37,
    input logic [DATA_WIDTH-1:0] data38,
    input logic [DATA_WIDTH-1:0] data39,
    input logic [DATA_WIDTH-1:0] data40,
    input logic [DATA_WIDTH-1:0] data41,
    input logic [DATA_WIDTH-1:0] data42,
    input logic [DATA_WIDTH-1:0] data43,
    input logic [DATA_WIDTH-1:0] data44,
    input logic [DATA_WIDTH-1:0] data45,
    input logic [DATA_WIDTH-1:0] data46,
    input logic [DATA_WIDTH-1:0] data47,
    input logic [DATA_WIDTH-1:0] data48,
    input logic [DATA_WIDTH-1:0] data49,
    input logic [DATA_WIDTH-1:0] data50,
    input logic [DATA_WIDTH-1:0] data51,
    input logic [DATA_WIDTH-1:0] data52,
    input logic [DATA_WIDTH-1:0] data53,
    input logic [DATA_WIDTH-1:0] data54,
    input logic [DATA_WIDTH-1:0] data55,
    input logic [DATA_WIDTH-1:0] data56,
    input logic [DATA_WIDTH-1:0] data57,
    input logic [DATA_WIDTH-1:0] data58,
    input logic [DATA_WIDTH-1:0] data59,
    input logic [DATA_WIDTH-1:0] data60,
    input logic [DATA_WIDTH-1:0] data61,
    input logic [DATA_WIDTH-1:0] data62,
    input logic [DATA_WIDTH-1:0] data63,
    input valid_in,
    input clk,
    input rst_n,
    output reg [31:0] data_out_1,
    output reg [31:0] data_out_2,
    output reg [31:0] data_out_3,
    output reg [31:0] data_out_4,
    output reg [31:0] data_out_5,
    output reg [31:0] data_out_6,
    output reg [31:0] data_out_7,
    output reg [31:0] data_out_8,
    output reg [31:0] data_out_9,
    output reg [31:0] data_out_10,
    output reg [31:0] data_out_11,
    output reg [31:0] data_out_12,
    output reg [31:0] data_out_13,
    output reg [31:0] data_out_14,
    output reg [31:0] data_out_15,
    output reg [31:0] data_out_16,
    output reg [31:0] data_out_17,
    output reg [31:0] data_out_18,
    output reg [31:0] data_out_19,
    output reg [31:0] data_out_20,
    output reg [31:0] data_out_21,
    output reg [31:0] data_out_22,
    output reg [31:0] data_out_23,
    output reg [31:0] data_out_24,
    output reg [31:0] data_out_25,
    output reg [31:0] data_out_26,
    output reg [31:0] data_out_27,
    output reg [31:0] data_out_28,
    output reg [31:0] data_out_29,
    output reg [31:0] data_out_30,
    output reg [31:0] data_out_31,
    output reg [31:0] data_out_32,
    output reg [31:0] data_out_33,
    output reg [31:0] data_out_34,
    output reg [31:0] data_out_35,
    output reg [31:0] data_out_36,
    output reg [31:0] data_out_37,
    output reg [31:0] data_out_38,
    output reg [31:0] data_out_39,
    output reg [31:0] data_out_40,
    output reg [31:0] data_out_41,
    output reg [31:0] data_out_42,
    output reg [31:0] data_out_43,
    output reg [31:0] data_out_44,
    output reg [31:0] data_out_45,
    output reg [31:0] data_out_46,
    output reg [31:0] data_out_47,
    output reg [31:0] data_out_48,
    output reg [31:0] data_out_49,
    output reg [31:0] data_out_50,
    output reg [31:0] data_out_51,
    output reg [31:0] data_out_52,
    output reg [31:0] data_out_53,
    output reg [31:0] data_out_54,
    output reg [31:0] data_out_55,
    output reg [31:0] data_out_56,
    output reg [31:0] data_out_57,
    output reg [31:0] data_out_58,
    output reg [31:0] data_out_59,
    output reg [31:0] data_out_60,
    output reg [31:0] data_out_61,
    output reg [31:0] data_out_62,
    output reg [31:0] data_out_63,
    output reg [31:0] data_out_64,
    output reg [31:0] data_out_65,
    output reg [31:0] data_out_66,
    output reg [31:0] data_out_67,
    output reg [31:0] data_out_68,
    output reg [31:0] data_out_69,
    output reg [31:0] data_out_70,
    output reg [31:0] data_out_71,
    output reg [31:0] data_out_72,
    output reg [31:0] data_out_73,
    output reg [31:0] data_out_74,
    output reg [31:0] data_out_75,
    output reg [31:0] data_out_76,
    output reg [31:0] data_out_77,
    output reg [31:0] data_out_78,
    output reg [31:0] data_out_79,
    output reg [31:0] data_out_80,
    output reg [31:0] data_out_81,
    output reg [31:0] data_out_82,
    output reg [31:0] data_out_83,
    output reg [31:0] data_out_84,
    output reg [31:0] data_out_85,
    output reg [31:0] data_out_86,
    output reg [31:0] data_out_87,
    output reg [31:0] data_out_88,
    output reg [31:0] data_out_89,
    output reg [31:0] data_out_90,
    output reg [31:0] data_out_91,
    output reg [31:0] data_out_92,
    output reg [31:0] data_out_93,
    output reg [31:0] data_out_94,
    output reg [31:0] data_out_95,
    output reg [31:0] data_out_96,
    output reg [31:0] data_out_97,
    output reg [31:0] data_out_98,
    output reg [31:0] data_out_99,
    output reg [31:0] data_out_100,
    output reg [31:0] data_out_101,
    output reg [31:0] data_out_102,
    output reg [31:0] data_out_103,
    output reg [31:0] data_out_104,
    output reg [31:0] data_out_105,
    output reg [31:0] data_out_106,
    output reg [31:0] data_out_107,
    output reg [31:0] data_out_108,
    output reg [31:0] data_out_109,
    output reg [31:0] data_out_110,
    output reg [31:0] data_out_111,
    output reg [31:0] data_out_112,
    output reg [31:0] data_out_113,
    output reg [31:0] data_out_114,
    output reg [31:0] data_out_115,
    output reg [31:0] data_out_116,
    output reg [31:0] data_out_117,
    output reg [31:0] data_out_118,
    output reg [31:0] data_out_119,
    output reg [31:0] data_out_120,
    output reg [31:0] data_out_121,
    output reg [31:0] data_out_122,
    output reg [31:0] data_out_123,
    output reg [31:0] data_out_124,
    output reg [31:0] data_out_125,
    output reg [31:0] data_out_126,
    output reg [31:0] data_out_127,
    output reg [31:0] data_out_128,          
    output reg valid_out_layer3
    
    );
    
    
reg valid_out_input_buffer;
 reg [31:0] buffer0 [0:7][0:5];  // 채널 0의 버퍼
    reg [31:0] buffer1 [0:7][0:5];  // 채널 1의 버퍼
    reg [31:0] buffer2 [0:7][0:5];  // 채널 2의 버퍼
    reg [31:0] buffer3 [0:7][0:5];  // 채널 3의 버퍼
    reg [31:0] buffer4 [0:7][0:5];  // 채널 4의 버퍼
    reg [31:0] buffer5 [0:7][0:5];  // 채널 5의 버퍼
    reg [31:0] buffer6 [0:7][0:5];  // 채널 6의 버퍼
    reg [31:0] buffer7 [0:7][0:5];  // 채널 7의 버퍼
    reg [31:0] buffer8 [0:7][0:5];  // 채널 8의 버퍼
    reg [31:0] buffer9 [0:7][0:5];  // 채널 9의 버퍼
    reg [31:0] buffer10 [0:7][0:5]; // 채널 10의 버퍼
    reg [31:0] buffer11 [0:7][0:5]; // 채널 11의 버퍼
    reg [31:0] buffer12 [0:7][0:5]; // 채널 12의 버퍼
    reg [31:0] buffer13 [0:7][0:5]; // 채널 13의 버퍼
    reg [31:0] buffer14 [0:7][0:5]; // 채널 14의 버퍼
    reg [31:0] buffer15 [0:7][0:5]; // 채널 15의 버퍼
    reg [31:0] buffer16 [0:7][0:5]; // 채널 16의 버퍼
    reg [31:0] buffer17 [0:7][0:5]; // 채널 17의 버퍼
    reg [31:0] buffer18 [0:7][0:5]; // 채널 18의 버퍼
    reg [31:0] buffer19 [0:7][0:5]; // 채널 19의 버퍼
    reg [31:0] buffer20 [0:7][0:5]; // 채널 20의 버퍼
    reg [31:0] buffer21 [0:7][0:5]; // 채널 21의 버퍼
    reg [31:0] buffer22 [0:7][0:5]; // 채널 22의 버퍼
    reg [31:0] buffer23 [0:7][0:5]; // 채널 23의 버퍼
    reg [31:0] buffer24 [0:7][0:5]; // 채널 24의 버퍼
    reg [31:0] buffer25 [0:7][0:5]; // 채널 25의 버퍼
    reg [31:0] buffer26 [0:7][0:5]; // 채널 26의 버퍼
    reg [31:0] buffer27 [0:7][0:5]; // 채널 27의 버퍼
    reg [31:0] buffer28 [0:7][0:5]; // 채널 28의 버퍼
    reg [31:0] buffer29 [0:7][0:5]; // 채널 29의 버퍼
    reg [31:0] buffer30 [0:7][0:5]; // 채널 30의 버퍼
    reg [31:0] buffer31 [0:7][0:5]; // 채널 31의 버퍼    
    reg [31:0] buffer32 [0:7][0:5]; // 채널 24의 버퍼
    reg [31:0] buffer33 [0:7][0:5]; // 채널 25의 버퍼
    reg [31:0] buffer34 [0:7][0:5]; // 채널 26의 버퍼
    reg [31:0] buffer35 [0:7][0:5]; // 채널 27의 버퍼
    reg [31:0] buffer36 [0:7][0:5]; // 채널 28의 버퍼
    reg [31:0] buffer37 [0:7][0:5]; // 채널 29의 버퍼
    reg [31:0] buffer38 [0:7][0:5]; // 채널 30의 버퍼
    reg [31:0] buffer39 [0:7][0:5]; // 채널 31의 버퍼  
    reg [31:0] buffer40 [0:7][0:5]; // 채널 24의 버퍼
    reg [31:0] buffer41 [0:7][0:5]; // 채널 25의 버퍼
    reg [31:0] buffer42 [0:7][0:5]; // 채널 26의 버퍼
    reg [31:0] buffer43 [0:7][0:5]; // 채널 27의 버퍼
    reg [31:0] buffer44 [0:7][0:5]; // 채널 28의 버퍼
    reg [31:0] buffer45 [0:7][0:5]; // 채널 29의 버퍼
    reg [31:0] buffer46 [0:7][0:5]; // 채널 30의 버퍼
    reg [31:0] buffer47 [0:7][0:5]; // 채널 31의 버퍼  
    reg [31:0] buffer48 [0:7][0:5]; // 채널 24의 버퍼
    reg [31:0] buffer49 [0:7][0:5]; // 채널 25의 버퍼
    reg [31:0] buffer50 [0:7][0:5]; // 채널 26의 버퍼
    reg [31:0] buffer51 [0:7][0:5]; // 채널 27의 버퍼
    reg [31:0] buffer52 [0:7][0:5]; // 채널 28의 버퍼
    reg [31:0] buffer53 [0:7][0:5]; // 채널 29의 버퍼
    reg [31:0] buffer54 [0:7][0:5]; // 채널 30의 버퍼
    reg [31:0] buffer55 [0:7][0:5]; // 채널 31의 버퍼  
    reg [31:0] buffer56 [0:7][0:5]; // 채널 24의 버퍼
    reg [31:0] buffer57 [0:7][0:5]; // 채널 25의 버퍼
    reg [31:0] buffer58 [0:7][0:5]; // 채널 26의 버퍼
    reg [31:0] buffer59 [0:7][0:5]; // 채널 27의 버퍼
    reg [31:0] buffer60 [0:7][0:5]; // 채널 28의 버퍼
    reg [31:0] buffer61 [0:7][0:5]; // 채널 29의 버퍼
    reg [31:0] buffer62 [0:7][0:5]; // 채널 30의 버퍼
    reg [31:0] buffer63 [0:7][0:5]; // 채널 31의 버퍼  
    
    reg valid_out_zero_padding_third;
    reg [31:0] padded0  [0:9][0:7];  // 패딩 0
    reg [31:0] padded1  [0:9][0:7];  // 패딩 1
    reg [31:0] padded2  [0:9][0:7];  // 패딩 2
    reg [31:0] padded3  [0:9][0:7];  // 패딩 3
    reg [31:0] padded4  [0:9][0:7];  // 패딩 4
    reg [31:0] padded5  [0:9][0:7];  // 패딩 5
    reg [31:0] padded6  [0:9][0:7];  // 패딩 6
    reg [31:0] padded7  [0:9][0:7];  // 패딩 7
    reg [31:0] padded8  [0:9][0:7];  // 패딩 8
    reg [31:0] padded9  [0:9][0:7];  // 패딩 9
    reg [31:0] padded10 [0:9][0:7];  // 패딩 10
    reg [31:0] padded11 [0:9][0:7];  // 패딩 11
    reg [31:0] padded12 [0:9][0:7];  // 패딩 12
    reg [31:0] padded13 [0:9][0:7];  // 패딩 13
    reg [31:0] padded14 [0:9][0:7];  // 패딩 14
    reg [31:0] padded15 [0:9][0:7];  // 패딩 15
    reg [31:0] padded16 [0:9][0:7];  // 패딩 16
    reg [31:0] padded17 [0:9][0:7];  // 패딩 17
    reg [31:0] padded18 [0:9][0:7];  // 패딩 18
    reg [31:0] padded19 [0:9][0:7];  // 패딩 19
    reg [31:0] padded20 [0:9][0:7];  // 패딩 20
    reg [31:0] padded21 [0:9][0:7];  // 패딩 21
    reg [31:0] padded22 [0:9][0:7];  // 패딩 22
    reg [31:0] padded23 [0:9][0:7];  // 패딩 23
    reg [31:0] padded24 [0:9][0:7];  // 패딩 24
    reg [31:0] padded25 [0:9][0:7];  // 패딩 25
    reg [31:0] padded26 [0:9][0:7];  // 패딩 26
    reg [31:0] padded27 [0:9][0:7];  // 패딩 27
    reg [31:0] padded28 [0:9][0:7];  // 패딩 28
    reg [31:0] padded29 [0:9][0:7];  // 패딩 29
    reg [31:0] padded30 [0:9][0:7];  // 패딩 30
    reg [31:0] padded31 [0:9][0:7];  // 패딩 31
    reg [31:0] padded32 [0:9][0:7];  // 패딩 1
    reg [31:0] padded33 [0:9][0:7];  // 패딩 2
    reg [31:0] padded34  [0:9][0:7];  // 패딩 3
    reg [31:0] padded35  [0:9][0:7];  // 패딩 4
    reg [31:0] padded36  [0:9][0:7];  // 패딩 5
    reg [31:0] padded37 [0:9][0:7];  // 패딩 6
    reg [31:0] padded38 [0:9][0:7];  // 패딩 7
    reg [31:0] padded39  [0:9][0:7];  // 패딩 8
    reg [31:0] padded40  [0:9][0:7];  // 패딩 9
    reg [31:0] padded41 [0:9][0:7];  // 패딩 10
    reg [31:0] padded42 [0:9][0:7];  // 패딩 11
    reg [31:0] padded43 [0:9][0:7];  // 패딩 12
    reg [31:0] padded44 [0:9][0:7];  // 패딩 13
    reg [31:0] padded45 [0:9][0:7];  // 패딩 14
    reg [31:0] padded46 [0:9][0:7];  // 패딩 15
    reg [31:0] padded47 [0:9][0:7];  // 패딩 16
    reg [31:0] padded48 [0:9][0:7];  // 패딩 17
    reg [31:0] padded49 [0:9][0:7];  // 패딩 18
    reg [31:0] padded50 [0:9][0:7];  // 패딩 19
    reg [31:0] padded51 [0:9][0:7];  // 패딩 20
    reg [31:0] padded52 [0:9][0:7];  // 패딩 21
    reg [31:0] padded53 [0:9][0:7];  // 패딩 22
    reg [31:0] padded54 [0:9][0:7];  // 패딩 23
    reg [31:0] padded55 [0:9][0:7];  // 패딩 24
    reg [31:0] padded56 [0:9][0:7];  // 패딩 25
    reg [31:0] padded57 [0:9][0:7];  // 패딩 26
    reg [31:0] padded58 [0:9][0:7];  // 패딩 27
    reg [31:0] padded59 [0:9][0:7];  // 패딩 28
    reg [31:0] padded60 [0:9][0:7];  // 패딩 29
    reg [31:0] padded61 [0:9][0:7];  // 패딩 30
    reg [31:0] padded62 [0:9][0:7];  // 패딩 31
    reg [31:0] padded63  [0:9][0:7];  // 패딩 0
    reg valid_out_threebythree;
    reg [DATA_WIDTH-1:0] patch [0:2][0:2];
    
    reg [31:0] data_out_conv3 [0:127];
    reg valid_out_conv3;
    
    reg [31:0] data_out_conv3_accum [0:127];
    reg valid_out_conv3_accum;
    
    reg [31:0] data_out_relu3 [0:127];
    reg valid_out_relu3;    
    
    reg [31:0] data_out_buf_1  [0:1][0:1];
reg [31:0] data_out_buf_2  [0:1][0:1];
reg [31:0] data_out_buf_3  [0:1][0:1];
reg [31:0] data_out_buf_4  [0:1][0:1];
reg [31:0] data_out_buf_5  [0:1][0:1];
reg [31:0] data_out_buf_6  [0:1][0:1];
reg [31:0] data_out_buf_7  [0:1][0:1];
reg [31:0] data_out_buf_8  [0:1][0:1];
reg [31:0] data_out_buf_9  [0:1][0:1];
reg [31:0] data_out_buf_10 [0:1][0:1];
reg [31:0] data_out_buf_11 [0:1][0:1];
reg [31:0] data_out_buf_12 [0:1][0:1];
reg [31:0] data_out_buf_13 [0:1][0:1];
reg [31:0] data_out_buf_14 [0:1][0:1];
reg [31:0] data_out_buf_15 [0:1][0:1];
reg [31:0] data_out_buf_16 [0:1][0:1];
reg [31:0] data_out_buf_17 [0:1][0:1];
reg [31:0] data_out_buf_18 [0:1][0:1];
reg [31:0] data_out_buf_19 [0:1][0:1];
reg [31:0] data_out_buf_20 [0:1][0:1];
reg [31:0] data_out_buf_21 [0:1][0:1];
reg [31:0] data_out_buf_22 [0:1][0:1];
reg [31:0] data_out_buf_23 [0:1][0:1];
reg [31:0] data_out_buf_24 [0:1][0:1];
reg [31:0] data_out_buf_25 [0:1][0:1];
reg [31:0] data_out_buf_26 [0:1][0:1];
reg [31:0] data_out_buf_27 [0:1][0:1];
reg [31:0] data_out_buf_28 [0:1][0:1];
reg [31:0] data_out_buf_29 [0:1][0:1];
reg [31:0] data_out_buf_30 [0:1][0:1];
reg [31:0] data_out_buf_31 [0:1][0:1];
reg [31:0] data_out_buf_32 [0:1][0:1];
reg [31:0] data_out_buf_33 [0:1][0:1];
reg [31:0] data_out_buf_34 [0:1][0:1];
reg [31:0] data_out_buf_35 [0:1][0:1];
reg [31:0] data_out_buf_36 [0:1][0:1];
reg [31:0] data_out_buf_37 [0:1][0:1];
reg [31:0] data_out_buf_38 [0:1][0:1];
reg [31:0] data_out_buf_39 [0:1][0:1];
reg [31:0] data_out_buf_40 [0:1][0:1];
reg [31:0] data_out_buf_41 [0:1][0:1];
reg [31:0] data_out_buf_42 [0:1][0:1];
reg [31:0] data_out_buf_43 [0:1][0:1];
reg [31:0] data_out_buf_44 [0:1][0:1];
reg [31:0] data_out_buf_45 [0:1][0:1];
reg [31:0] data_out_buf_46 [0:1][0:1];
reg [31:0] data_out_buf_47 [0:1][0:1];
reg [31:0] data_out_buf_48 [0:1][0:1];
reg [31:0] data_out_buf_49 [0:1][0:1];
reg [31:0] data_out_buf_50 [0:1][0:1];
reg [31:0] data_out_buf_51 [0:1][0:1];
reg [31:0] data_out_buf_52 [0:1][0:1];
reg [31:0] data_out_buf_53 [0:1][0:1];
reg [31:0] data_out_buf_54 [0:1][0:1];
reg [31:0] data_out_buf_55 [0:1][0:1];
reg [31:0] data_out_buf_56 [0:1][0:1];
reg [31:0] data_out_buf_57 [0:1][0:1];
reg [31:0] data_out_buf_58 [0:1][0:1];
reg [31:0] data_out_buf_59 [0:1][0:1];
reg [31:0] data_out_buf_60 [0:1][0:1];
reg [31:0] data_out_buf_61 [0:1][0:1];
reg [31:0] data_out_buf_62 [0:1][0:1];
reg [31:0] data_out_buf_63 [0:1][0:1];
reg [31:0] data_out_buf_64 [0:1][0:1];
reg [31:0] data_out_buf_65 [0:1][0:1];
reg [31:0] data_out_buf_66 [0:1][0:1];
reg [31:0] data_out_buf_67 [0:1][0:1];
reg [31:0] data_out_buf_68 [0:1][0:1];
reg [31:0] data_out_buf_69 [0:1][0:1];
reg [31:0] data_out_buf_70 [0:1][0:1];
reg [31:0] data_out_buf_71 [0:1][0:1];
reg [31:0] data_out_buf_72 [0:1][0:1];
reg [31:0] data_out_buf_73 [0:1][0:1];
reg [31:0] data_out_buf_74 [0:1][0:1];
reg [31:0] data_out_buf_75 [0:1][0:1];
reg [31:0] data_out_buf_76 [0:1][0:1];
reg [31:0] data_out_buf_77 [0:1][0:1];
reg [31:0] data_out_buf_78 [0:1][0:1];
reg [31:0] data_out_buf_79 [0:1][0:1];
reg [31:0] data_out_buf_80 [0:1][0:1];
reg [31:0] data_out_buf_81 [0:1][0:1];
reg [31:0] data_out_buf_82 [0:1][0:1];
reg [31:0] data_out_buf_83 [0:1][0:1];
reg [31:0] data_out_buf_84 [0:1][0:1];
reg [31:0] data_out_buf_85 [0:1][0:1];
reg [31:0] data_out_buf_86 [0:1][0:1];
reg [31:0] data_out_buf_87 [0:1][0:1];
reg [31:0] data_out_buf_88 [0:1][0:1];
reg [31:0] data_out_buf_89 [0:1][0:1];
reg [31:0] data_out_buf_90 [0:1][0:1];
reg [31:0] data_out_buf_91 [0:1][0:1];
reg [31:0] data_out_buf_92 [0:1][0:1];
reg [31:0] data_out_buf_93 [0:1][0:1];
reg [31:0] data_out_buf_94 [0:1][0:1];
reg [31:0] data_out_buf_95 [0:1][0:1];
reg [31:0] data_out_buf_96 [0:1][0:1];
reg [31:0] data_out_buf_97 [0:1][0:1];
reg [31:0] data_out_buf_98 [0:1][0:1];
reg [31:0] data_out_buf_99 [0:1][0:1];
reg [31:0] data_out_buf_100 [0:1][0:1];
reg [31:0] data_out_buf_101 [0:1][0:1];
reg [31:0] data_out_buf_102 [0:1][0:1];
reg [31:0] data_out_buf_103 [0:1][0:1];
reg [31:0] data_out_buf_104 [0:1][0:1];
reg [31:0] data_out_buf_105 [0:1][0:1];
reg [31:0] data_out_buf_106 [0:1][0:1];
reg [31:0] data_out_buf_107 [0:1][0:1];
reg [31:0] data_out_buf_108 [0:1][0:1];
reg [31:0] data_out_buf_109 [0:1][0:1];
reg [31:0] data_out_buf_110 [0:1][0:1];
reg [31:0] data_out_buf_111 [0:1][0:1];
reg [31:0] data_out_buf_112 [0:1][0:1];
reg [31:0] data_out_buf_113 [0:1][0:1];
reg [31:0] data_out_buf_114 [0:1][0:1];
reg [31:0] data_out_buf_115 [0:1][0:1];
reg [31:0] data_out_buf_116 [0:1][0:1];
reg [31:0] data_out_buf_117 [0:1][0:1];
reg [31:0] data_out_buf_118 [0:1][0:1];
reg [31:0] data_out_buf_119 [0:1][0:1];
reg [31:0] data_out_buf_120 [0:1][0:1];
reg [31:0] data_out_buf_121 [0:1][0:1];
reg [31:0] data_out_buf_122 [0:1][0:1];
reg [31:0] data_out_buf_123 [0:1][0:1];
reg [31:0] data_out_buf_124 [0:1][0:1];
reg [31:0] data_out_buf_125 [0:1][0:1];
reg [31:0] data_out_buf_126 [0:1][0:1];
reg [31:0] data_out_buf_127 [0:1][0:1];
reg [31:0] data_out_buf_128 [0:1][0:1];
reg valid_out_channel_buffer3;

input_buffer_3 #(
.DATA_WIDTH(32),
.CHANNELS(64),
.WIDTH(6),
.HEIGHT(8)
)input_buffer_3(
.valid_in(valid_in),
.data0(data0),
.data1(data1),
.data2(data2),
.data3(data3),
.data4(data4),
.data5(data5),
.data6(data6),
.data7(data7),
.data8(data8),
.data9(data9),
.data10(data10),
.data11(data11),
.data12(data12),
.data13(data13),
.data14(data14),
.data15(data15),
.data16(data16),
.data17(data17),
.data18(data18),
.data19(data19),
.data20(data20),
.data21(data21),
.data22(data22),
.data23(data23),
.data24(data24),
.data25(data25),
.data26(data26),
.data27(data27),
.data28(data28),
.data29(data29),
.data30(data30),
.data31(data31),
.data32(data32),
.data33(data33),
.data34(data34),
.data35(data35),
.data36(data36),
.data37(data37),
.data38(data38),
.data39(data39),
.data40(data40),
.data41(data41),
.data42(data42),
.data43(data43),
.data44(data44),
.data45(data45),
.data46(data46),
.data47(data47),
.data48(data48),
.data49(data49),
.data50(data50),
.data51(data51),
.data52(data52),
.data53(data53),
.data54(data54),
.data55(data55),
.data56(data56),
.data57(data57),
.data58(data58),
.data59(data59),
.data60(data60),
.data61(data61),
.data62(data62),
.data63(data63),
.clk(clk),
.rst_n(rst_n),
.buffer0(buffer0),
.buffer1(buffer1),
.buffer2(buffer2),
.buffer3(buffer3),
.buffer4(buffer4),
.buffer5(buffer5),
.buffer6(buffer6),
.buffer7(buffer7),
.buffer8(buffer8),
.buffer9(buffer9),
.buffer10(buffer10),
.buffer11(buffer11),
.buffer12(buffer12),
.buffer13(buffer13),
.buffer14(buffer14),
.buffer15(buffer15),
.buffer16(buffer16),
.buffer17(buffer17),
.buffer18(buffer18),
.buffer19(buffer19),
.buffer20(buffer20),
.buffer21(buffer21),
.buffer22(buffer22),
.buffer23(buffer23),
.buffer24(buffer24),
.buffer25(buffer25),
.buffer26(buffer26),
.buffer27(buffer27),
.buffer28(buffer28),
.buffer29(buffer29),
.buffer30(buffer30),
.buffer31(buffer31),
.buffer32(buffer32),
.buffer33(buffer33),
.buffer34(buffer34),
.buffer35(buffer35),
.buffer36(buffer36),
.buffer37(buffer37),
.buffer38(buffer38),
.buffer39(buffer39),
.buffer40(buffer40),
.buffer41(buffer41),
.buffer42(buffer42),
.buffer43(buffer43),
.buffer44(buffer44),
.buffer45(buffer45),
.buffer46(buffer46),
.buffer47(buffer47),
.buffer48(buffer48),
.buffer49(buffer49),
.buffer50(buffer50),
.buffer51(buffer51),
.buffer52(buffer52),
.buffer53(buffer53),
.buffer54(buffer54),
.buffer55(buffer55),
.buffer56(buffer56),
.buffer57(buffer57),
.buffer58(buffer58),
.buffer59(buffer59),
.buffer60(buffer60),
.buffer61(buffer61),
.buffer62(buffer62),
.buffer63(buffer63),
.valid_out(valid_out_input_buffer)
);

zero_padding_third #(
.DATA_WIDTH(32),
.PAD_WIDTH(8),
.PAD_HEIGHT(10),
.WIDTH(6),
.HEIGHT(8)
)zero_padding_third(
 .buffer0(buffer0),
.buffer1(buffer1),
.buffer2(buffer2),
.buffer3(buffer3),
.buffer4(buffer4),
.buffer5(buffer5),
.buffer6(buffer6),
.buffer7(buffer7),
.buffer8(buffer8),
.buffer9(buffer9),
.buffer10(buffer10),
.buffer11(buffer11),
.buffer12(buffer12),
.buffer13(buffer13),
.buffer14(buffer14),
.buffer15(buffer15),
.buffer16(buffer16),
.buffer17(buffer17),
.buffer18(buffer18),
.buffer19(buffer19),
.buffer20(buffer20),
.buffer21(buffer21),
.buffer22(buffer22),
.buffer23(buffer23),
.buffer24(buffer24),
.buffer25(buffer25),
.buffer26(buffer26),
.buffer27(buffer27),
.buffer28(buffer28),
.buffer29(buffer29),
.buffer30(buffer30),
.buffer31(buffer31),
.buffer32(buffer32),
.buffer33(buffer33),
.buffer34(buffer34),
.buffer35(buffer35),
.buffer36(buffer36),
.buffer37(buffer37),
.buffer38(buffer38),
.buffer39(buffer39),
.buffer40(buffer40),
.buffer41(buffer41),
.buffer42(buffer42),
.buffer43(buffer43),
.buffer44(buffer44),
.buffer45(buffer45),
.buffer46(buffer46),
.buffer47(buffer47),
.buffer48(buffer48),
.buffer49(buffer49),
.buffer50(buffer50),
.buffer51(buffer51),
.buffer52(buffer52),
.buffer53(buffer53),
.buffer54(buffer54),
.buffer55(buffer55),
.buffer56(buffer56),
.buffer57(buffer57),
.buffer58(buffer58),
.buffer59(buffer59),
.buffer60(buffer60),
.buffer61(buffer61),
.buffer62(buffer62),
.buffer63(buffer63),
.valid_in(valid_out_input_buffer),
.rst_n(rst_n),
.clk(clk),
.padded0(padded0),
.padded1(padded1),
.padded2(padded2),
.padded3(padded3),
.padded4(padded4),
.padded5(padded5),
.padded6(padded6),
.padded7(padded7),
.padded8(padded8),
.padded9(padded9),
.padded10(padded10),
.padded11(padded11),
.padded12(padded12),
.padded13(padded13),
.padded14(padded14),
.padded15(padded15),
.padded16(padded16),
.padded17(padded17),
.padded18(padded18),
.padded19(padded19),
.padded20(padded20),
.padded21(padded21),
.padded22(padded22),
.padded23(padded23),
.padded24(padded24),
.padded25(padded25),
.padded26(padded26),
.padded27(padded27),
.padded28(padded28),
.padded29(padded29),
.padded30(padded30),
.padded31(padded31),
.padded32(padded32),
.padded33(padded33),
.padded34(padded34),
.padded35(padded35),
.padded36(padded36),
.padded37(padded37),
.padded38(padded38),
.padded39(padded39),
.padded40(padded40),
.padded41(padded41),
.padded42(padded42),
.padded43(padded43),
.padded44(padded44),
.padded45(padded45),
.padded46(padded46),
.padded47(padded47),
.padded48(padded48),
.padded49(padded49),
.padded50(padded50),
.padded51(padded51),
.padded52(padded52),
.padded53(padded53),
.padded54(padded54),
.padded55(padded55),
.padded56(padded56),
.padded57(padded57),
.padded58(padded58),
.padded59(padded59),
.padded60(padded60),
.padded61(padded61),
.padded62(padded62),
.padded63(padded63),
.valid_padding(valid_out_zero_padding_third)
);

threebythree_3 #(
.DATA_WIDTH(32),
.PAD_WIDTH(8),
.PAD_HEIGHT(10)
)threebythree_3(
.padded0(padded0),
.padded1(padded1),
.padded2(padded2),
.padded3(padded3),
.padded4(padded4),
.padded5(padded5),
.padded6(padded6),
.padded7(padded7),
.padded8(padded8),
.padded9(padded9),
.padded10(padded10),
.padded11(padded11),
.padded12(padded12),
.padded13(padded13),
.padded14(padded14),
.padded15(padded15),
.padded16(padded16),
.padded17(padded17),
.padded18(padded18),
.padded19(padded19),
.padded20(padded20),
.padded21(padded21),
.padded22(padded22),
.padded23(padded23),
.padded24(padded24),
.padded25(padded25),
.padded26(padded26),
.padded27(padded27),
.padded28(padded28),
.padded29(padded29),
.padded30(padded30),
.padded31(padded31),
.padded32(padded32),
.padded33(padded33),
.padded34(padded34),
.padded35(padded35),
.padded36(padded36),
.padded37(padded37),
.padded38(padded38),
.padded39(padded39),
.padded40(padded40),
.padded41(padded41),
.padded42(padded42),
.padded43(padded43),
.padded44(padded44),
.padded45(padded45),
.padded46(padded46),
.padded47(padded47),
.padded48(padded48),
.padded49(padded49),
.padded50(padded50),
.padded51(padded51),
.padded52(padded52),
.padded53(padded53),
.padded54(padded54),
.padded55(padded55),
.padded56(padded56),
.padded57(padded57),
.padded58(padded58),
.padded59(padded59),
.padded60(padded60),
.padded61(padded61),
.padded62(padded62),
.padded63(padded63),
.valid_padding(valid_out_zero_padding_third),
.rst_n(rst_n),
.clk(clk),
.patch(patch),
.valid_out(valid_out_threebythree)
);

conv3_layer conv3_layer(
.clk(clk),
.rst_n(rst_n),
.valid_in(valid_out_threebythree),
.data_in(patch),
.conv3_out(data_out_conv3),
.valid_out(valid_out_conv3)
);

conv3_accum #(
.WIDTH(6),
.HEIGHT(8),
.SIZE(48),
.filter_num(128),
.channel_num(64)
) conv3_accum(
.data_in(data_out_conv3),
.valid_in(valid_out_conv3),
.clk(clk),
.rst_n(rst_n),
.data_out(data_out_conv3_accum),
.valid_out(valid_out_conv3_accum)
);

relu3#(
.IMAGE_WIDTH(6),
.IMAGE_HEIGHT(8),
.CHANNELS(128),
.DATA_BITS(32)
)relu3(
.data_in(data_out_conv3_accum),
.valid_in(valid_out_conv3_accum),
.rst_n(rst_n),
.clk(clk),
.data_out(data_out_relu3),
.valid_out(valid_out_relu3)
);

channel_buffer3#(
.IMAGE_WIDTH(6),
.IMAGE_HEIGHT(8),
.CHANNELS(128),
.DATA_BITS(32)
)channel_buffer3(
.data_in(data_out_relu3),
.valid_in(valid_out_relu3),
.clk(clk),
.rst_n(rst_n),
.data_out_1(data_out_buf_1),
.data_out_2(data_out_buf_2),
.data_out_3(data_out_buf_3),
.data_out_4(data_out_buf_4),
.data_out_5(data_out_buf_5),
.data_out_6(data_out_buf_6),
.data_out_7(data_out_buf_7),
.data_out_8(data_out_buf_8),
.data_out_9(data_out_buf_9),
.data_out_10(data_out_buf_10),
.data_out_11(data_out_buf_11),
.data_out_12(data_out_buf_12),
.data_out_13(data_out_buf_13),
.data_out_14(data_out_buf_14),
.data_out_15(data_out_buf_15),
.data_out_16(data_out_buf_16),
.data_out_17(data_out_buf_17),
.data_out_18(data_out_buf_18),
.data_out_19(data_out_buf_19),
.data_out_20(data_out_buf_20),
.data_out_21(data_out_buf_21),
.data_out_22(data_out_buf_22),
.data_out_23(data_out_buf_23),
.data_out_24(data_out_buf_24),
.data_out_25(data_out_buf_25),
.data_out_26(data_out_buf_26),
.data_out_27(data_out_buf_27),
.data_out_28(data_out_buf_28),
.data_out_29(data_out_buf_29),
.data_out_30(data_out_buf_30),
.data_out_31(data_out_buf_31),
.data_out_32(data_out_buf_32),
.data_out_33(data_out_buf_33),
.data_out_34(data_out_buf_34),
.data_out_35(data_out_buf_35),
.data_out_36(data_out_buf_36),
.data_out_37(data_out_buf_37),
.data_out_38(data_out_buf_38),
.data_out_39(data_out_buf_39),
.data_out_40(data_out_buf_40),
.data_out_41(data_out_buf_41),
.data_out_42(data_out_buf_42),
.data_out_43(data_out_buf_43),
.data_out_44(data_out_buf_44),
.data_out_45(data_out_buf_45),
.data_out_46(data_out_buf_46),
.data_out_47(data_out_buf_47),
.data_out_48(data_out_buf_48),
.data_out_49(data_out_buf_49),
.data_out_50(data_out_buf_50),
.data_out_51(data_out_buf_51),
.data_out_52(data_out_buf_52),
.data_out_53(data_out_buf_53),
.data_out_54(data_out_buf_54),
.data_out_55(data_out_buf_55),
.data_out_56(data_out_buf_56),
.data_out_57(data_out_buf_57),
.data_out_58(data_out_buf_58),
.data_out_59(data_out_buf_59),
.data_out_60(data_out_buf_60),
.data_out_61(data_out_buf_61),
.data_out_62(data_out_buf_62),
.data_out_63(data_out_buf_63),
.data_out_64(data_out_buf_64),
.data_out_65(data_out_buf_65),
.data_out_66(data_out_buf_66),
.data_out_67(data_out_buf_67),
.data_out_68(data_out_buf_68),
.data_out_69(data_out_buf_69),
.data_out_70(data_out_buf_70),
.data_out_71(data_out_buf_71),
.data_out_72(data_out_buf_72),
.data_out_73(data_out_buf_73),
.data_out_74(data_out_buf_74),
.data_out_75(data_out_buf_75),
.data_out_76(data_out_buf_76),
.data_out_77(data_out_buf_77),
.data_out_78(data_out_buf_78),
.data_out_79(data_out_buf_79),
.data_out_80(data_out_buf_80),
.data_out_81(data_out_buf_81),
.data_out_82(data_out_buf_82),
.data_out_83(data_out_buf_83),
.data_out_84(data_out_buf_84),
.data_out_85(data_out_buf_85),
.data_out_86(data_out_buf_86),
.data_out_87(data_out_buf_87),
.data_out_88(data_out_buf_88),
.data_out_89(data_out_buf_89),
.data_out_90(data_out_buf_90),
.data_out_91(data_out_buf_91),
.data_out_92(data_out_buf_92),
.data_out_93(data_out_buf_93),
.data_out_94(data_out_buf_94),
.data_out_95(data_out_buf_95),
.data_out_96(data_out_buf_96),
.data_out_97(data_out_buf_97),
.data_out_98(data_out_buf_98),
.data_out_99(data_out_buf_99),
.data_out_100(data_out_buf_100),
.data_out_101(data_out_buf_101),
.data_out_102(data_out_buf_102),
.data_out_103(data_out_buf_103),
.data_out_104(data_out_buf_104),
.data_out_105(data_out_buf_105),
.data_out_106(data_out_buf_106),
.data_out_107(data_out_buf_107),
.data_out_108(data_out_buf_108),
.data_out_109(data_out_buf_109),
.data_out_110(data_out_buf_110),
.data_out_111(data_out_buf_111),
.data_out_112(data_out_buf_112),
.data_out_113(data_out_buf_113),
.data_out_114(data_out_buf_114),
.data_out_115(data_out_buf_115),
.data_out_116(data_out_buf_116),
.data_out_117(data_out_buf_117),
.data_out_118(data_out_buf_118),
.data_out_119(data_out_buf_119),
.data_out_120(data_out_buf_120),
.data_out_121(data_out_buf_121),
.data_out_122(data_out_buf_122),
.data_out_123(data_out_buf_123),
.data_out_124(data_out_buf_124),
.data_out_125(data_out_buf_125),
.data_out_126(data_out_buf_126),
.data_out_127(data_out_buf_127),
.data_out_128(data_out_buf_128),
.valid_out(valid_out_channel_buffer3)
);

max_pooling_layer_top3 max_pooling_layer_top3(
.valid_in(valid_out_channel_buffer3),
.rst_n(rst_n),
.clk(clk),
.valid_out(valid_out_layer3),
.data_in_1(data_out_buf_1),
.data_in_2(data_out_buf_2),
.data_in_3(data_out_buf_3),
.data_in_4(data_out_buf_4),
.data_in_5(data_out_buf_5),
.data_in_6(data_out_buf_6),
.data_in_7(data_out_buf_7),
.data_in_8(data_out_buf_8),
.data_in_9(data_out_buf_9),
.data_in_10(data_out_buf_10),
.data_in_11(data_out_buf_11),
.data_in_12(data_out_buf_12),
.data_in_13(data_out_buf_13),
.data_in_14(data_out_buf_14),
.data_in_15(data_out_buf_15),
.data_in_16(data_out_buf_16),
.data_in_17(data_out_buf_17),
.data_in_18(data_out_buf_18),
.data_in_19(data_out_buf_19),
.data_in_20(data_out_buf_20),
.data_in_21(data_out_buf_21),
.data_in_22(data_out_buf_22),
.data_in_23(data_out_buf_23),
.data_in_24(data_out_buf_24),
.data_in_25(data_out_buf_25),
.data_in_26(data_out_buf_26),
.data_in_27(data_out_buf_27),
.data_in_28(data_out_buf_28),
.data_in_29(data_out_buf_29),
.data_in_30(data_out_buf_30),
.data_in_31(data_out_buf_31),
.data_in_32(data_out_buf_32),
.data_in_33(data_out_buf_33),
.data_in_34(data_out_buf_34),
.data_in_35(data_out_buf_35),
.data_in_36(data_out_buf_36),
.data_in_37(data_out_buf_37),
.data_in_38(data_out_buf_38),
.data_in_39(data_out_buf_39),
.data_in_40(data_out_buf_40),
.data_in_41(data_out_buf_41),
.data_in_42(data_out_buf_42),
.data_in_43(data_out_buf_43),
.data_in_44(data_out_buf_44),
.data_in_45(data_out_buf_45),
.data_in_46(data_out_buf_46),
.data_in_47(data_out_buf_47),
.data_in_48(data_out_buf_48),
.data_in_49(data_out_buf_49),
.data_in_50(data_out_buf_50),
.data_in_51(data_out_buf_51),
.data_in_52(data_out_buf_52),
.data_in_53(data_out_buf_53),
.data_in_54(data_out_buf_54),
.data_in_55(data_out_buf_55),
.data_in_56(data_out_buf_56),
.data_in_57(data_out_buf_57),
.data_in_58(data_out_buf_58),
.data_in_59(data_out_buf_59),
.data_in_60(data_out_buf_60),
.data_in_61(data_out_buf_61),
.data_in_62(data_out_buf_62),
.data_in_63(data_out_buf_63),
.data_in_64(data_out_buf_64),
.data_in_65(data_out_buf_65),
.data_in_66(data_out_buf_66),
.data_in_67(data_out_buf_67),
.data_in_68(data_out_buf_68),
.data_in_69(data_out_buf_69),
.data_in_70(data_out_buf_70),
.data_in_71(data_out_buf_71),
.data_in_72(data_out_buf_72),
.data_in_73(data_out_buf_73),
.data_in_74(data_out_buf_74),
.data_in_75(data_out_buf_75),
.data_in_76(data_out_buf_76),
.data_in_77(data_out_buf_77),
.data_in_78(data_out_buf_78),
.data_in_79(data_out_buf_79),
.data_in_80(data_out_buf_80),
.data_in_81(data_out_buf_81),
.data_in_82(data_out_buf_82),
.data_in_83(data_out_buf_83),
.data_in_84(data_out_buf_84),
.data_in_85(data_out_buf_85),
.data_in_86(data_out_buf_86),
.data_in_87(data_out_buf_87),
.data_in_88(data_out_buf_88),
.data_in_89(data_out_buf_89),
.data_in_90(data_out_buf_90),
.data_in_91(data_out_buf_91),
.data_in_92(data_out_buf_92),
.data_in_93(data_out_buf_93),
.data_in_94(data_out_buf_94),
.data_in_95(data_out_buf_95),
.data_in_96(data_out_buf_96),
.data_in_97(data_out_buf_97),
.data_in_98(data_out_buf_98),
.data_in_99(data_out_buf_99),
.data_in_100(data_out_buf_100),
.data_in_101(data_out_buf_101),
.data_in_102(data_out_buf_102),
.data_in_103(data_out_buf_103),
.data_in_104(data_out_buf_104),
.data_in_105(data_out_buf_105),
.data_in_106(data_out_buf_106),
.data_in_107(data_out_buf_107),
.data_in_108(data_out_buf_108),
.data_in_109(data_out_buf_109),
.data_in_110(data_out_buf_110),
.data_in_111(data_out_buf_111),
.data_in_112(data_out_buf_112),
.data_in_113(data_out_buf_113),
.data_in_114(data_out_buf_114),
.data_in_115(data_out_buf_115),
.data_in_116(data_out_buf_116),
.data_in_117(data_out_buf_117),
.data_in_118(data_out_buf_118),
.data_in_119(data_out_buf_119),
.data_in_120(data_out_buf_120),
.data_in_121(data_out_buf_121),
.data_in_122(data_out_buf_122),
.data_in_123(data_out_buf_123),
.data_in_124(data_out_buf_124),
.data_in_125(data_out_buf_125),
.data_in_126(data_out_buf_126),
.data_in_127(data_out_buf_127),
.data_in_128(data_out_buf_128),
.data_out_1(data_out_1),
.data_out_2(data_out_2),
.data_out_3(data_out_3),
.data_out_4(data_out_4),
.data_out_5(data_out_5),
.data_out_6(data_out_6),
.data_out_7(data_out_7),
.data_out_8(data_out_8),
.data_out_9(data_out_9),
.data_out_10(data_out_10),
.data_out_11(data_out_11),
.data_out_12(data_out_12),
.data_out_13(data_out_13),
.data_out_14(data_out_14),
.data_out_15(data_out_15),
.data_out_16(data_out_16),
.data_out_17(data_out_17),
.data_out_18(data_out_18),
.data_out_19(data_out_19),
.data_out_20(data_out_20),
.data_out_21(data_out_21),
.data_out_22(data_out_22),
.data_out_23(data_out_23),
.data_out_24(data_out_24),
.data_out_25(data_out_25),
.data_out_26(data_out_26),
.data_out_27(data_out_27),
.data_out_28(data_out_28),
.data_out_29(data_out_29),
.data_out_30(data_out_30),
.data_out_31(data_out_31),
.data_out_32(data_out_32),
.data_out_33(data_out_33),
.data_out_34(data_out_34),
.data_out_35(data_out_35),
.data_out_36(data_out_36),
.data_out_37(data_out_37),
.data_out_38(data_out_38),
.data_out_39(data_out_39),
.data_out_40(data_out_40),
.data_out_41(data_out_41),
.data_out_42(data_out_42),
.data_out_43(data_out_43),
.data_out_44(data_out_44),
.data_out_45(data_out_45),
.data_out_46(data_out_46),
.data_out_47(data_out_47),
.data_out_48(data_out_48),
.data_out_49(data_out_49),
.data_out_50(data_out_50),
.data_out_51(data_out_51),
.data_out_52(data_out_52),
.data_out_53(data_out_53),
.data_out_54(data_out_54),
.data_out_55(data_out_55),
.data_out_56(data_out_56),
.data_out_57(data_out_57),
.data_out_58(data_out_58),
.data_out_59(data_out_59),
.data_out_60(data_out_60),
.data_out_61(data_out_61),
.data_out_62(data_out_62),
.data_out_63(data_out_63),
.data_out_64(data_out_64),
.data_out_65(data_out_65),
.data_out_66(data_out_66),
.data_out_67(data_out_67),
.data_out_68(data_out_68),
.data_out_69(data_out_69),
.data_out_70(data_out_70),
.data_out_71(data_out_71),
.data_out_72(data_out_72),
.data_out_73(data_out_73),
.data_out_74(data_out_74),
.data_out_75(data_out_75),
.data_out_76(data_out_76),
.data_out_77(data_out_77),
.data_out_78(data_out_78),
.data_out_79(data_out_79),
.data_out_80(data_out_80),
.data_out_81(data_out_81),
.data_out_82(data_out_82),
.data_out_83(data_out_83),
.data_out_84(data_out_84),
.data_out_85(data_out_85),
.data_out_86(data_out_86),
.data_out_87(data_out_87),
.data_out_88(data_out_88),
.data_out_89(data_out_89),
.data_out_90(data_out_90),
.data_out_91(data_out_91),
.data_out_92(data_out_92),
.data_out_93(data_out_93),
.data_out_94(data_out_94),
.data_out_95(data_out_95),
.data_out_96(data_out_96),
.data_out_97(data_out_97),
.data_out_98(data_out_98),
.data_out_99(data_out_99),
.data_out_100(data_out_100),
.data_out_101(data_out_101),
.data_out_102(data_out_102),
.data_out_103(data_out_103),
.data_out_104(data_out_104),
.data_out_105(data_out_105),
.data_out_106(data_out_106),
.data_out_107(data_out_107),
.data_out_108(data_out_108),
.data_out_109(data_out_109),
.data_out_110(data_out_110),
.data_out_111(data_out_111),
.data_out_112(data_out_112),
.data_out_113(data_out_113),
.data_out_114(data_out_114),
.data_out_115(data_out_115),
.data_out_116(data_out_116),
.data_out_117(data_out_117),
.data_out_118(data_out_118),
.data_out_119(data_out_119),
.data_out_120(data_out_120),
.data_out_121(data_out_121),
.data_out_122(data_out_122),
.data_out_123(data_out_123),
.data_out_124(data_out_124),
.data_out_125(data_out_125),
.data_out_126(data_out_126),
.data_out_127(data_out_127),
.data_out_128(data_out_128)
);

endmodule
