`timescale 1ns / 1ps

module max_pooling_layer_top3 (
    input wire clk,
    input wire rst_n,
    input wire valid_in,
    input wire [31:0] data_in_1 [0:1][0:1],
    input wire [31:0] data_in_2 [0:1][0:1],
    input wire [31:0] data_in_3 [0:1][0:1],
    input wire [31:0] data_in_4 [0:1][0:1],
    input wire [31:0] data_in_5 [0:1][0:1],
    input wire [31:0] data_in_6 [0:1][0:1],
    input wire [31:0] data_in_7 [0:1][0:1],
    input wire [31:0] data_in_8 [0:1][0:1],
    input wire [31:0] data_in_9 [0:1][0:1],
    input wire [31:0] data_in_10 [0:1][0:1],
    input wire [31:0] data_in_11 [0:1][0:1],
    input wire [31:0] data_in_12 [0:1][0:1],
    input wire [31:0] data_in_13 [0:1][0:1],
    input wire [31:0] data_in_14 [0:1][0:1],
    input wire [31:0] data_in_15 [0:1][0:1],
    input wire [31:0] data_in_16 [0:1][0:1],
    input wire [31:0] data_in_17 [0:1][0:1],
    input wire [31:0] data_in_18 [0:1][0:1],
    input wire [31:0] data_in_19 [0:1][0:1],
    input wire [31:0] data_in_20 [0:1][0:1],
    input wire [31:0] data_in_21 [0:1][0:1],
    input wire [31:0] data_in_22 [0:1][0:1],
    input wire [31:0] data_in_23 [0:1][0:1],
    input wire [31:0] data_in_24 [0:1][0:1],
    input wire [31:0] data_in_25 [0:1][0:1],
    input wire [31:0] data_in_26 [0:1][0:1],
    input wire [31:0] data_in_27 [0:1][0:1],
    input wire [31:0] data_in_28 [0:1][0:1],
    input wire [31:0] data_in_29 [0:1][0:1],
    input wire [31:0] data_in_30 [0:1][0:1],
    input wire [31:0] data_in_31 [0:1][0:1],
    input wire [31:0] data_in_32 [0:1][0:1],
    input wire [31:0] data_in_33 [0:1][0:1],
    input wire [31:0] data_in_34 [0:1][0:1],
    input wire [31:0] data_in_35 [0:1][0:1],
    input wire [31:0] data_in_36 [0:1][0:1],
    input wire [31:0] data_in_37 [0:1][0:1],
    input wire [31:0] data_in_38 [0:1][0:1],
    input wire [31:0] data_in_39 [0:1][0:1],
    input wire [31:0] data_in_40 [0:1][0:1],
    input wire [31:0] data_in_41 [0:1][0:1],
    input wire [31:0] data_in_42 [0:1][0:1],
    input wire [31:0] data_in_43 [0:1][0:1],
    input wire [31:0] data_in_44 [0:1][0:1],
    input wire [31:0] data_in_45 [0:1][0:1],
    input wire [31:0] data_in_46 [0:1][0:1],
    input wire [31:0] data_in_47 [0:1][0:1],
    input wire [31:0] data_in_48 [0:1][0:1],
    input wire [31:0] data_in_49 [0:1][0:1],
    input wire [31:0] data_in_50 [0:1][0:1],
    input wire [31:0] data_in_51 [0:1][0:1],
    input wire [31:0] data_in_52 [0:1][0:1],
    input wire [31:0] data_in_53 [0:1][0:1],
    input wire [31:0] data_in_54 [0:1][0:1],
    input wire [31:0] data_in_55 [0:1][0:1],
    input wire [31:0] data_in_56 [0:1][0:1],
    input wire [31:0] data_in_57 [0:1][0:1],
    input wire [31:0] data_in_58 [0:1][0:1],
    input wire [31:0] data_in_59 [0:1][0:1],
    input wire [31:0] data_in_60 [0:1][0:1],
    input wire [31:0] data_in_61 [0:1][0:1],
    input wire [31:0] data_in_62 [0:1][0:1],
    input wire [31:0] data_in_63 [0:1][0:1],
    input wire [31:0] data_in_64 [0:1][0:1],
    input wire [31:0] data_in_65 [0:1][0:1],
input wire [31:0] data_in_66 [0:1][0:1],
input wire [31:0] data_in_67 [0:1][0:1],
input wire [31:0] data_in_68 [0:1][0:1],
input wire [31:0] data_in_69 [0:1][0:1],
input wire [31:0] data_in_70 [0:1][0:1],
input wire [31:0] data_in_71 [0:1][0:1],
input wire [31:0] data_in_72 [0:1][0:1],
input wire [31:0] data_in_73 [0:1][0:1],
input wire [31:0] data_in_74 [0:1][0:1],
input wire [31:0] data_in_75 [0:1][0:1],
input wire [31:0] data_in_76 [0:1][0:1],
input wire [31:0] data_in_77 [0:1][0:1],
input wire [31:0] data_in_78 [0:1][0:1],
input wire [31:0] data_in_79 [0:1][0:1],
input wire [31:0] data_in_80 [0:1][0:1],
input wire [31:0] data_in_81 [0:1][0:1],
input wire [31:0] data_in_82 [0:1][0:1],
input wire [31:0] data_in_83 [0:1][0:1],
input wire [31:0] data_in_84 [0:1][0:1],
input wire [31:0] data_in_85 [0:1][0:1],
input wire [31:0] data_in_86 [0:1][0:1],
input wire [31:0] data_in_87 [0:1][0:1],
input wire [31:0] data_in_88 [0:1][0:1],
input wire [31:0] data_in_89 [0:1][0:1],
input wire [31:0] data_in_90 [0:1][0:1],
input wire [31:0] data_in_91 [0:1][0:1],
input wire [31:0] data_in_92 [0:1][0:1],
input wire [31:0] data_in_93 [0:1][0:1],
input wire [31:0] data_in_94 [0:1][0:1],
input wire [31:0] data_in_95 [0:1][0:1],
input wire [31:0] data_in_96 [0:1][0:1],
input wire [31:0] data_in_97 [0:1][0:1],
input wire [31:0] data_in_98 [0:1][0:1],
input wire [31:0] data_in_99 [0:1][0:1],
input wire [31:0] data_in_100 [0:1][0:1],
input wire [31:0] data_in_101 [0:1][0:1],
input wire [31:0] data_in_102 [0:1][0:1],
input wire [31:0] data_in_103 [0:1][0:1],
input wire [31:0] data_in_104 [0:1][0:1],
input wire [31:0] data_in_105 [0:1][0:1],
input wire [31:0] data_in_106 [0:1][0:1],
input wire [31:0] data_in_107 [0:1][0:1],
input wire [31:0] data_in_108 [0:1][0:1],
input wire [31:0] data_in_109 [0:1][0:1],
input wire [31:0] data_in_110 [0:1][0:1],
input wire [31:0] data_in_111 [0:1][0:1],
input wire [31:0] data_in_112 [0:1][0:1],
input wire [31:0] data_in_113 [0:1][0:1],
input wire [31:0] data_in_114 [0:1][0:1],
input wire [31:0] data_in_115 [0:1][0:1],
input wire [31:0] data_in_116 [0:1][0:1],
input wire [31:0] data_in_117 [0:1][0:1],
input wire [31:0] data_in_118 [0:1][0:1],
input wire [31:0] data_in_119 [0:1][0:1],
input wire [31:0] data_in_120 [0:1][0:1],
input wire [31:0] data_in_121 [0:1][0:1],
input wire [31:0] data_in_122 [0:1][0:1],
input wire [31:0] data_in_123 [0:1][0:1],
input wire [31:0] data_in_124 [0:1][0:1],
input wire [31:0] data_in_125 [0:1][0:1],
input wire [31:0] data_in_126 [0:1][0:1],
input wire [31:0] data_in_127 [0:1][0:1],
input wire [31:0] data_in_128 [0:1][0:1],
    output reg [31:0] data_out_1,
    output reg [31:0] data_out_2,
    output reg [31:0] data_out_3,
    output reg [31:0] data_out_4,
    output reg [31:0] data_out_5,
    output reg [31:0] data_out_6,
    output reg [31:0] data_out_7,
    output reg [31:0] data_out_8,
    output reg [31:0] data_out_9,
    output reg [31:0] data_out_10,
    output reg [31:0] data_out_11,
    output reg [31:0] data_out_12,
    output reg [31:0] data_out_13,
    output reg [31:0] data_out_14,
    output reg [31:0] data_out_15,
    output reg [31:0] data_out_16,
    output reg [31:0] data_out_17,
    output reg [31:0] data_out_18,
    output reg [31:0] data_out_19,
    output reg [31:0] data_out_20,
    output reg [31:0] data_out_21,
    output reg [31:0] data_out_22,
    output reg [31:0] data_out_23,
    output reg [31:0] data_out_24,
    output reg [31:0] data_out_25,
    output reg [31:0] data_out_26,
    output reg [31:0] data_out_27,
    output reg [31:0] data_out_28,
    output reg [31:0] data_out_29,
    output reg [31:0] data_out_30,
    output reg [31:0] data_out_31,
    output reg [31:0] data_out_32,
    output reg [31:0] data_out_33,
    output reg [31:0] data_out_34,
    output reg [31:0] data_out_35,
    output reg [31:0] data_out_36,
    output reg [31:0] data_out_37,
    output reg [31:0] data_out_38,
    output reg [31:0] data_out_39,
    output reg [31:0] data_out_40,
    output reg [31:0] data_out_41,
    output reg [31:0] data_out_42,
    output reg [31:0] data_out_43,
    output reg [31:0] data_out_44,
    output reg [31:0] data_out_45,
    output reg [31:0] data_out_46,
    output reg [31:0] data_out_47,
    output reg [31:0] data_out_48,
    output reg [31:0] data_out_49,
    output reg [31:0] data_out_50,
    output reg [31:0] data_out_51,
    output reg [31:0] data_out_52,
    output reg [31:0] data_out_53,
    output reg [31:0] data_out_54,
    output reg [31:0] data_out_55,
    output reg [31:0] data_out_56,
    output reg [31:0] data_out_57,
    output reg [31:0] data_out_58,
    output reg [31:0] data_out_59,
    output reg [31:0] data_out_60,
    output reg [31:0] data_out_61,
    output reg [31:0] data_out_62,
    output reg [31:0] data_out_63,
    output reg [31:0] data_out_64,
    output reg [31:0] data_out_65,
output reg [31:0] data_out_66,
output reg [31:0] data_out_67,
output reg [31:0] data_out_68,
output reg [31:0] data_out_69,
output reg [31:0] data_out_70,
output reg [31:0] data_out_71,
output reg [31:0] data_out_72,
output reg [31:0] data_out_73,
output reg [31:0] data_out_74,
output reg [31:0] data_out_75,
output reg [31:0] data_out_76,
output reg [31:0] data_out_77,
output reg [31:0] data_out_78,
output reg [31:0] data_out_79,
output reg [31:0] data_out_80,
output reg [31:0] data_out_81,
output reg [31:0] data_out_82,
output reg [31:0] data_out_83,
output reg [31:0] data_out_84,
output reg [31:0] data_out_85,
output reg [31:0] data_out_86,
output reg [31:0] data_out_87,
output reg [31:0] data_out_88,
output reg [31:0] data_out_89,
output reg [31:0] data_out_90,
output reg [31:0] data_out_91,
output reg [31:0] data_out_92,
output reg [31:0] data_out_93,
output reg [31:0] data_out_94,
output reg [31:0] data_out_95,
output reg [31:0] data_out_96,
output reg [31:0] data_out_97,
output reg [31:0] data_out_98,
output reg [31:0] data_out_99,
output reg [31:0] data_out_100,
output reg [31:0] data_out_101,
output reg [31:0] data_out_102,
output reg [31:0] data_out_103,
output reg [31:0] data_out_104,
output reg [31:0] data_out_105,
output reg [31:0] data_out_106,
output reg [31:0] data_out_107,
output reg [31:0] data_out_108,
output reg [31:0] data_out_109,
output reg [31:0] data_out_110,
output reg [31:0] data_out_111,
output reg [31:0] data_out_112,
output reg [31:0] data_out_113,
output reg [31:0] data_out_114,
output reg [31:0] data_out_115,
output reg [31:0] data_out_116,
output reg [31:0] data_out_117,
output reg [31:0] data_out_118,
output reg [31:0] data_out_119,
output reg [31:0] data_out_120,
output reg [31:0] data_out_121,
output reg [31:0] data_out_122,
output reg [31:0] data_out_123,
output reg [31:0] data_out_124,
output reg [31:0] data_out_125,
output reg [31:0] data_out_126,
output reg [31:0] data_out_127,
output reg [31:0] data_out_128,
    output reg valid_out
);
integer delay;
reg cnt[1:0];
    // 각 max_pooling 모듈에 들어가는 입력을 설정하는 블록
    reg [31:0] data_in_i [0:127][0:1][0:1];

    // 각 max_pooling 모듈에서 나오는 출력
    reg [31:0] max_out [0:127];

    // Generate 블록에서 각 입력 값을 설정
    generate
        genvar i;
        for (i = 0; i < 128; i = i + 1) begin : gen_max_pooling
            always @(*) begin
            if(valid_in == 1) begin
                case(i)
                    0: data_in_i[i] = data_in_1;
                    1: data_in_i[i] = data_in_2;
                    2: data_in_i[i] = data_in_3;
                    3: data_in_i[i] = data_in_4;
                    4: data_in_i[i] = data_in_5;
                    5: data_in_i[i] = data_in_6;
                    6: data_in_i[i] = data_in_7;
                    7: data_in_i[i] = data_in_8;
                    8: data_in_i[i] = data_in_9;
                    9: data_in_i[i] = data_in_10;
                    10: data_in_i[i] = data_in_11;
                    11: data_in_i[i] = data_in_12;
                    12: data_in_i[i] = data_in_13;
                    13: data_in_i[i] = data_in_14;
                    14: data_in_i[i] = data_in_15;
                    15: data_in_i[i] = data_in_16;
                    16: data_in_i[i] = data_in_17;
                    17: data_in_i[i] = data_in_18;
                    18: data_in_i[i] = data_in_19;
                    19: data_in_i[i] = data_in_20;
                    20: data_in_i[i] = data_in_21;
                    21: data_in_i[i] = data_in_22;
                    22: data_in_i[i] = data_in_23;
                    23: data_in_i[i] = data_in_24;
                    24: data_in_i[i] = data_in_25;
                    25: data_in_i[i] = data_in_26;
                    26: data_in_i[i] = data_in_27;
                    27: data_in_i[i] = data_in_28;
                    28: data_in_i[i] = data_in_29;
                    29: data_in_i[i] = data_in_30;
                    30: data_in_i[i] = data_in_31;
                    31: data_in_i[i] = data_in_32;
                    32: data_in_i[i] = data_in_33;
                    33: data_in_i[i] = data_in_34;
                    34: data_in_i[i] = data_in_35;
                    35: data_in_i[i] = data_in_36;
                    36: data_in_i[i] = data_in_37;
                    37: data_in_i[i] = data_in_38;
                    38: data_in_i[i] = data_in_39;
                    39: data_in_i[i] = data_in_40;
                    40: data_in_i[i] = data_in_41;
                    41: data_in_i[i] = data_in_42;
                    42: data_in_i[i] = data_in_43;
                    43: data_in_i[i] = data_in_44;
                    44: data_in_i[i] = data_in_45;
                    45: data_in_i[i] = data_in_46;
                    46: data_in_i[i] = data_in_47;
                    47: data_in_i[i] = data_in_48;
                    48: data_in_i[i] = data_in_49;
                    49: data_in_i[i] = data_in_50;
                    50: data_in_i[i] = data_in_51;
                    51: data_in_i[i] = data_in_52;
                    52: data_in_i[i] = data_in_53;
                    53: data_in_i[i] = data_in_54;
                    54: data_in_i[i] = data_in_55;
                    55: data_in_i[i] = data_in_56;
                    56: data_in_i[i] = data_in_57;
                    57: data_in_i[i] = data_in_58;
                    58: data_in_i[i] = data_in_59;
                    59: data_in_i[i] = data_in_60;
                    60: data_in_i[i] = data_in_61;
                    61: data_in_i[i] = data_in_62;
                    62: data_in_i[i] = data_in_63;
                    63: data_in_i[i] = data_in_64;
                    64: data_in_i[i] = data_in_65;
                    65: data_in_i[i] = data_in_66;
                    66: data_in_i[i] = data_in_67;
                    67: data_in_i[i] = data_in_68;
                    68: data_in_i[i] = data_in_69;
                    69: data_in_i[i] = data_in_70;
                    70: data_in_i[i] = data_in_71;
                    71: data_in_i[i] = data_in_72;
                    72: data_in_i[i] = data_in_73;
                    73: data_in_i[i] = data_in_74;
                    74: data_in_i[i] = data_in_75;
                    75: data_in_i[i] = data_in_76;
                    76: data_in_i[i] = data_in_77;
                    77: data_in_i[i] = data_in_78;
                    78: data_in_i[i] = data_in_79;
                    79: data_in_i[i] = data_in_80;
                    80: data_in_i[i] = data_in_81;
                    81: data_in_i[i] = data_in_82;
                    82: data_in_i[i] = data_in_83;
                    83: data_in_i[i] = data_in_84;
                    84: data_in_i[i] = data_in_85;
                    85: data_in_i[i] = data_in_86;
                    86: data_in_i[i] = data_in_87;
                    87: data_in_i[i] = data_in_88;
                    88: data_in_i[i] = data_in_89;
                    89: data_in_i[i] = data_in_90;
                    90: data_in_i[i] = data_in_91;
                    91: data_in_i[i] = data_in_92;
                    92: data_in_i[i] = data_in_93;
                    93: data_in_i[i] = data_in_94;                                                 
                    94: data_in_i[i] = data_in_95;
                    95: data_in_i[i] = data_in_96;
                    96: data_in_i[i] = data_in_97;
                    97: data_in_i[i] = data_in_98;
                    98: data_in_i[i] = data_in_99;
                    99: data_in_i[i] = data_in_100;
                    100: data_in_i[i] = data_in_101;
                    101: data_in_i[i] = data_in_102;
                    102: data_in_i[i] = data_in_103;
                    103: data_in_i[i] = data_in_104;
                    104: data_in_i[i] = data_in_105;
                    105: data_in_i[i] = data_in_106;
                    106: data_in_i[i] = data_in_107;
                    107: data_in_i[i] = data_in_108;
                    108: data_in_i[i] = data_in_109;
                    109: data_in_i[i] = data_in_110;
                    110: data_in_i[i] = data_in_111;
                    111: data_in_i[i] = data_in_112;
                    112: data_in_i[i] = data_in_113;
                    113: data_in_i[i] = data_in_114;
                    114: data_in_i[i] = data_in_115;
                    115: data_in_i[i] = data_in_116;
                    116: data_in_i[i] = data_in_117;
                    117: data_in_i[i] = data_in_118;
                    118: data_in_i[i] = data_in_119;
                    119: data_in_i[i] = data_in_120;
                    120: data_in_i[i] = data_in_121;
                    121: data_in_i[i] = data_in_122;
                    122: data_in_i[i] = data_in_123;
                    123: data_in_i[i] = data_in_124;
                    124: data_in_i[i] = data_in_125;
                    125: data_in_i[i] = data_in_126;
                    126: data_in_i[i] = data_in_127;
                    127: data_in_i[i] = data_in_128;                     
                endcase
                end
            end

            max_pooling u_max_pooling (
                .clk(clk),
                .rst_n(rst_n),
                .data_in0(data_in_i[i][0][0]),
                .data_in1(data_in_i[i][0][1]),
                .data_in2(data_in_i[i][1][0]),
                .data_in3(data_in_i[i][1][1]),
                .data_out(max_out[i])
            );
        end
    endgenerate

    // 출력 처리 블록
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            // Reset output
            data_out_1 <= 32'b0;
            data_out_2 <= 32'b0;
            data_out_3 <= 32'b0;
            data_out_4 <= 32'b0;
            data_out_5 <= 32'b0;
            data_out_6 <= 32'b0;
            data_out_7 <= 32'b0;
            data_out_8 <= 32'b0;
            data_out_9 <= 32'b0;
            data_out_10 <= 32'b0;
            data_out_11 <= 32'b0;
            data_out_12 <= 32'b0;
            data_out_13 <= 32'b0;
            data_out_14 <= 32'b0;
            data_out_15 <= 32'b0;
            data_out_16 <= 32'b0;
            data_out_17 <= 32'b0;
            data_out_18 <= 32'b0;
            data_out_19 <= 32'b0;
            data_out_20 <= 32'b0;
            data_out_21 <= 32'b0;
            data_out_22 <= 32'b0;
            data_out_23 <= 32'b0;
            data_out_24 <= 32'b0;
            data_out_25 <= 32'b0;
            data_out_26 <= 32'b0;
            data_out_27 <= 32'b0;
            data_out_28 <= 32'b0;
            data_out_29 <= 32'b0;
            data_out_30 <= 32'b0;
            data_out_31 <= 32'b0;
            data_out_32 <= 32'b0;
            data_out_33 <= 32'b0;
            data_out_34 <= 32'b0;
            data_out_35 <= 32'b0;
            data_out_36 <= 32'b0;
            data_out_37 <= 32'b0;
            data_out_38 <= 32'b0;
            data_out_39 <= 32'b0;
            data_out_40 <= 32'b0;
            data_out_41 <= 32'b0;
            data_out_42 <= 32'b0;
            data_out_43 <= 32'b0;
            data_out_44 <= 32'b0;
            data_out_45 <= 32'b0;
            data_out_46 <= 32'b0;
            data_out_47 <= 32'b0;
            data_out_48 <= 32'b0;
            data_out_49 <= 32'b0;
            data_out_50 <= 32'b0;
            data_out_51 <= 32'b0;
            data_out_52 <= 32'b0;
            data_out_53 <= 32'b0;
            data_out_54 <= 32'b0;
            data_out_55 <= 32'b0;
            data_out_56 <= 32'b0;
            data_out_57 <= 32'b0;
            data_out_58 <= 32'b0;
            data_out_59 <= 32'b0;
            data_out_60 <= 32'b0;
            data_out_61 <= 32'b0;
            data_out_62 <= 32'b0;
            data_out_63 <= 32'b0;
            data_out_64 <= 32'b0;       
            data_out_65 <= 32'b0;
data_out_66 <= 32'b0;
data_out_67 <= 32'b0;
data_out_68 <= 32'b0;
data_out_69 <= 32'b0;
data_out_70 <= 32'b0;
data_out_71 <= 32'b0;
data_out_72 <= 32'b0;
data_out_73 <= 32'b0;
data_out_74 <= 32'b0;
data_out_75 <= 32'b0;
data_out_76 <= 32'b0;
data_out_77 <= 32'b0;
data_out_78 <= 32'b0;
data_out_79 <= 32'b0;
data_out_80 <= 32'b0;
data_out_81 <= 32'b0;
data_out_82 <= 32'b0;
data_out_83 <= 32'b0;
data_out_84 <= 32'b0;
data_out_85 <= 32'b0;
data_out_86 <= 32'b0;
data_out_87 <= 32'b0;
data_out_88 <= 32'b0;
data_out_89 <= 32'b0;
data_out_90 <= 32'b0;
data_out_91 <= 32'b0;
data_out_92 <= 32'b0;
data_out_93 <= 32'b0;
data_out_94 <= 32'b0;
data_out_95 <= 32'b0;
data_out_96 <= 32'b0;
data_out_97 <= 32'b0;
data_out_98 <= 32'b0;
data_out_99 <= 32'b0;
data_out_100 <= 32'b0;
data_out_101 <= 32'b0;
data_out_102 <= 32'b0;
data_out_103 <= 32'b0;
data_out_104 <= 32'b0;
data_out_105 <= 32'b0;
data_out_106 <= 32'b0;
data_out_107 <= 32'b0;
data_out_108 <= 32'b0;
data_out_109 <= 32'b0;
data_out_110 <= 32'b0;
data_out_111 <= 32'b0;
data_out_112 <= 32'b0;
data_out_113 <= 32'b0;
data_out_114 <= 32'b0;
data_out_115 <= 32'b0;
data_out_116 <= 32'b0;
data_out_117 <= 32'b0;
data_out_118 <= 32'b0;
data_out_119 <= 32'b0;
data_out_120 <= 32'b0;
data_out_121 <= 32'b0;
data_out_122 <= 32'b0;
data_out_123 <= 32'b0;
data_out_124 <= 32'b0;
data_out_125 <= 32'b0;
data_out_126 <= 32'b0;
data_out_127 <= 32'b0;
data_out_128 <= 32'b0;     
            valid_out <= 1'b0;
            cnt[0] <= 0;
            cnt[1] <= 1;
            
        end else begin
            data_out_1 <= max_out[0];
            data_out_2 <= max_out[1];
            data_out_3 <= max_out[2];
            data_out_4 <= max_out[3];
            data_out_5 <= max_out[4];
            data_out_6 <= max_out[5];
            data_out_7 <= max_out[6];
            data_out_8 <= max_out[7];
            data_out_9 <= max_out[8];
            data_out_10 <= max_out[9];
            data_out_11 <= max_out[10];
            data_out_12 <= max_out[11];
            data_out_13 <= max_out[12];
            data_out_14 <= max_out[13];
            data_out_15 <= max_out[14];
            data_out_16 <= max_out[15];
            data_out_17 <= max_out[16];
            data_out_18 <= max_out[17];
            data_out_19 <= max_out[18];
            data_out_20 <= max_out[19];
            data_out_21 <= max_out[20];
            data_out_22 <= max_out[21];
            data_out_23 <= max_out[22];
            data_out_24 <= max_out[23];
            data_out_25 <= max_out[24];
            data_out_26 <= max_out[25];
            data_out_27 <= max_out[26];
            data_out_28 <= max_out[27];
            data_out_29 <= max_out[28];
            data_out_30 <= max_out[29];
            data_out_31 <= max_out[30];
            data_out_32 <= max_out[31];
            data_out_33 <= max_out[32];
            data_out_34 <= max_out[33];
            data_out_35 <= max_out[34];
            data_out_36 <= max_out[35];
            data_out_37 <= max_out[36];
            data_out_38 <= max_out[37];
            data_out_39 <= max_out[38];
            data_out_40 <= max_out[39];
            data_out_41 <= max_out[40];
            data_out_42 <= max_out[41];
            data_out_43 <= max_out[42];
            data_out_44 <= max_out[43];
            data_out_45 <= max_out[44];
            data_out_46 <= max_out[45];
            data_out_47 <= max_out[46];
            data_out_48 <= max_out[47];
            data_out_49 <= max_out[48];
            data_out_50 <= max_out[49];
            data_out_51 <= max_out[50];
            data_out_52 <= max_out[51];
            data_out_53 <= max_out[52];
            data_out_54 <= max_out[53];
            data_out_55 <= max_out[54];
            data_out_56 <= max_out[55];
            data_out_57 <= max_out[56];
            data_out_58 <= max_out[57];
            data_out_59 <= max_out[58];
            data_out_60 <= max_out[59];
            data_out_61 <= max_out[60];
            data_out_62 <= max_out[61];
            data_out_63 <= max_out[62];
            data_out_64 <= max_out[63];
            data_out_65 <= max_out[64];
data_out_66 <= max_out[65];
data_out_67 <= max_out[66];
data_out_68 <= max_out[67];
data_out_69 <= max_out[68];
data_out_70 <= max_out[69];
data_out_71 <= max_out[70];
data_out_72 <= max_out[71];
data_out_73 <= max_out[72];
data_out_74 <= max_out[73];
data_out_75 <= max_out[74];
data_out_76 <= max_out[75];
data_out_77 <= max_out[76];
data_out_78 <= max_out[77];
data_out_79 <= max_out[78];
data_out_80 <= max_out[79];
data_out_81 <= max_out[80];
data_out_82 <= max_out[81];
data_out_83 <= max_out[82];
data_out_84 <= max_out[83];
data_out_85 <= max_out[84];
data_out_86 <= max_out[85];
data_out_87 <= max_out[86];
data_out_88 <= max_out[87];
data_out_89 <= max_out[88];
data_out_90 <= max_out[89];
data_out_91 <= max_out[90];
data_out_92 <= max_out[91];
data_out_93 <= max_out[92];
data_out_94 <= max_out[93];
data_out_95 <= max_out[94];
data_out_96 <= max_out[95];
data_out_97 <= max_out[96];
data_out_98 <= max_out[97];
data_out_99 <= max_out[98];
data_out_100 <= max_out[99];
data_out_101 <= max_out[100];
data_out_102 <= max_out[101];
data_out_103 <= max_out[102];
data_out_104 <= max_out[103];
data_out_105 <= max_out[104];
data_out_106 <= max_out[105];
data_out_107 <= max_out[106];
data_out_108 <= max_out[107];
data_out_109 <= max_out[108];
data_out_110 <= max_out[109];
data_out_111 <= max_out[110];
data_out_112 <= max_out[111];
data_out_113 <= max_out[112];
data_out_114 <= max_out[113];
data_out_115 <= max_out[114];
data_out_116 <= max_out[115];
data_out_117 <= max_out[116];
data_out_118 <= max_out[117];
data_out_119 <= max_out[118];
data_out_120 <= max_out[119];
data_out_121 <= max_out[120];
data_out_122 <= max_out[121];
data_out_123 <= max_out[122];
data_out_124 <= max_out[123];
data_out_125 <= max_out[124];
data_out_126 <= max_out[125];
data_out_127 <= max_out[126];
data_out_128 <= max_out[127];            
            
        end
        cnt[0] <= valid_in;
        cnt[1] <= cnt[0];
        assign valid_out = cnt[1];
        
    end
endmodule